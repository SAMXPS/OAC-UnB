-- ****************************************** 
--  Circuito: Memória RISCV 32
--  Autor: Samuel James de Lima Barroso / 190019948
-- ******************************************

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use std.textio.all;

entity memoriaRV is
    port (
        clock   : in  std_logic;
        wren    : in  std_logic;
        address : in  std_logic_vector; -- std_logic_vector sem tamanho pode ser utilizado para designar um
        datain  : in  std_logic_vector; -- tamanho flexível de dados, definido conforme a instância da arquitetura.
        dataout : out std_logic_vector
    );
end entity memoriaRV;

architecture memoriaRV_arch of memoriaRV is
    type   ram_type is array (0 to (2**address'length)-1) of std_logic_vector(datain'range);

    impure function init_ram_hex return ram_type  is
        file     text_file   : text open read_mode is "ram_content_hex.txt";
        variable text_line   : line;
        variable ram_depth   : natural := (2**address'length);
        variable ram_content : ram_type;
        begin
            for i in 0 to ram_depth - 1 loop
                readline(text_file, text_line);
                hread(text_line, ram_content(i));
            end loop;
            return ram_content;
    end function;

    signal mem : ram_type := init_ram_hex;
    signal read_address : std_logic_vector(address'range);

    begin

        dataout <= mem(to_integer(unsigned(read_address)));

        Write: process(clock) begin
            if wren = '1' then
                mem(to_integer(unsigned(address))) <= datain;
            end if;
            read_address <= address;
        end process;
end memoriaRV_arch;